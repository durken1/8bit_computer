library ieee;
use ieee.std_logic_1164.all;

package data_types is
  
  type output_en is (none, regA_o, regB_o, regI_o, alu_o);

end package;